`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    21:06:20 01/11/2018 
// Design Name: 
// Module Name:    U_MCB_WR 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module U_MCB_WR(
	input clk, 
	input rst_n,
	input u_wr_cmd_done,	//The operation of wirte cmd is done 
	input u_wr_rdy,				//user write ready ,data can be written in to mcb
	
	output reg u_wr_cmd_en,	//user write mcb cmd enable
	output reg u_wr_en,			//user write data enable
	output reg [127:0] u_wr_data,	//user write data
	output reg [29:0] u_wr_addr,	//user write address
	output reg [6:0] u_wr_len			//user write data len
    );
   
  (* KEEP = "TRUE" *) wire [1:0] u_wr_s_r;
	(* KEEP = "TRUE" *) wire [3:0] u_wr_en_dly1;
	
	parameter WR_IDLE 	= 2'd0,
						WR_BEGIN 	=	2'd1,
						WR_WAIT 	= 2'd2;
						
	reg [6:0] u_wr_cnt; //user write count	
	reg [1:0] u_wr_s; //user write state
	
	//when mcb write fifo more than 2 data enable write data cmd
	always@(posedge clk)
	begin
		if(!rst_n)
			begin
				u_wr_cmd_en <= 1'b0;
			end
		else
			begin
				if(u_wr_cmd_done)
					u_wr_cmd_en <= 1'b0;		//clear mcb user write enable signal
				else if(u_wr_cnt == 40)		
					u_wr_cmd_en <= 1'b1;	//enable user mcb cmd signal
			end
	end 
	
	
	//д��������
	
	always@(posedge clk)
	begin
		if(!rst_n)
		begin
			u_wr_data <= 128'hAA_AA_AA_AA_AA_AA_AA_AA_AA_AA_AA_AA_AA_AA_AA_AA;
		end
		else begin
			if(u_wr_rdy)							//mcb fifo is valid
				u_wr_data <= ~u_wr_data; // count up data write to mcb fifo
			else if(~u_wr_en)
				u_wr_data <= 128'hAA_AA_AA_AA_AA_AA_AA_AA_AA_AA_AA_AA_AA_AA_AA_AA;
		end
	end
	
	
	//д������
	
	always@(posedge clk)
	begin
		if(!rst_n)
			u_wr_cnt <= 7'd0;
		else begin
			if(u_wr_rdy) u_wr_cnt <= u_wr_cnt + 1'b1;
			else if (u_wr_s == WR_IDLE) u_wr_cnt <= 7'b0; 
		end
	end
	
	reg [29:0] u_wr_addr_set;
	
	//д����״̬��
	
	always@(posedge clk)
	begin
		if(!rst_n)
		begin
			u_wr_len <= 7'd64;			//user write len
			u_wr_addr <= 29'd0;			//user write addr
			u_wr_en <= 1'b0;				//user write enable
			u_wr_s <= WR_IDLE;
		end
		else begin
			case(u_wr_s)
				WR_IDLE:
				begin
					u_wr_en <= 1'b0;
					if(u_wr_cmd_en == 1'b0)	//start new write
						u_wr_s <= WR_BEGIN;
					else
						u_wr_s <= u_wr_s;
				end
				
				WR_BEGIN:
				begin
					u_wr_en <= 1'b1;
					u_wr_addr <= u_wr_addr_set;
					u_wr_len <= 7'd64;
					u_wr_s <= WR_WAIT;
				end
				
				WR_WAIT:
				begin
					if(u_wr_cnt == (u_wr_len - 1))
					begin
						u_wr_s <= WR_IDLE;
						u_wr_en <= 1'b0;
					end
					else u_wr_s <= u_wr_s;
				end
				
				default : u_wr_s <= WR_IDLE;
				
			endcase

		end

	end
	
	//��ַ�ռ���ʼ��ַ����
	parameter ADDR_INC = 12'h400;
	parameter END_ADDR = 29'h10000000 - ADDR_INC;
	
	always @(posedge clk)
	begin
		if(~rst_n)
		begin
			u_wr_addr_set <= 29'd0;
		end
		else begin
		if(u_wr_cmd_done && (u_wr_addr_set < END_ADDR))
			u_wr_addr_set <= u_wr_addr_set +  ADDR_INC;
		else if(u_wr_addr_set == END_ADDR)
			u_wr_addr_set <= 29'd0;
			
			
		end
		
		
		
		
	end
	
	
	
	
	
	
	
	

endmodule
