module Serial_Port_Driver(
	clk,
	rst_n,
	uart_tx_o,
	uart_rx_i,
	
	);












endmodule
